***PMOS characteristics
 vg 1 0 dc -2
 vd 3 0 dc -2.5
 v1 3 2 dc 0
.model pmod pmos level=54 version=4.7
 m1 0 1 2 2 pmod w=100u l=10u
.dc vg 0.0 -10.0 -0.1 
.control
 run
 plot  i(v1) xlabel 'vg' ylabel 'id' title 'transfer characteristics' 
.endc
.end