***characteristics of CMOS
 vg 1 0 dc 5
 vd 2 0 dc 5
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
 m1 3 1 0 0 nmod w=100u l=10u
 m2 3 1 2 2 pmod w=100u l=10u
 .dc vg 0 5 0.1
.control
 run
 plot v(1) v(3)   
.endc
.end










