***Transient Analysis
vin 2 0 pulse(0 5 0 0 0 100ms 200ms)
vin 2 0 5.0
 r1 2 1 1.2k
 c1 1 0 0.1u
 l1 1 0 100m
.tran 0.2ms 1000ms
.control
 run
plot v(1) v(2)
.endc
.end