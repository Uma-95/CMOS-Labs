***DC Analysis
vin 1 0 5.0
 r1 1 2 6k
 c1 2 0 18u
.dc vin 0.0 5.0 0.1
.control
 run
 plot v(1) v(2)
.endc
.end