***lab5_3
.subckt inverter 1 2 3
M1 3 1 2 2 pmod w=100u l=10u
M2 3 1 0 0 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.model pmod pmos version=54 level=4.7
.ends

.subckt pass_or 1 2 3 4
M1 2 2 4 4 nmod w=100u l=10u
M2 1 3 4 4 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.ends

.subckt pass_and 1 2 3 4
M1 2 3 4 4 nmod w=100u l=10u
M2 1 2 4 4 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.ends

Va 11 0 dc 0V
Vb 12 0 dc 0V
Vc 13 0 pulse (0 5 0 0 0 10m 20m)
Vd 14 0 dc 5V
Ve 15 0 dc 5V
Vdd 2 0 dc 5V
Xb 12 2 16 inverter
Xc 13 2 17 inverter
Xd 14 2 18 inverter
Xde 21 2 22 inverter
Xab 11 12 16 19 pass_and
Xabc 19 13 17 20 pass_or
Xabc_d 20 21 22 23 pass_and
.tran 0.1m 200m
.control 
run
plot V(23) V(13) 

.endc
.end