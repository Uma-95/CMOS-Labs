***AC Analysis
vin 1 0 dc 0 ac 5
 r1 1 2 8k
 r2 2 0 2k
.ac dec 10 1 10k
.control
 run
 plot v(1) v(2)
.endc
.end