
***ABC+D
.subckt inverter 1 2 3
M1 3 1 2 2 nmod w=100u l=10u
M2 3 1 0 0 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.model pmod pmos version=54 level=4.7
.ends

.subckt pass_or 1 2 3 4
M1 2 2 4 4 nmod w=100u l=10u
M2 1 3 4 4 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.ends

.subckt pass_and 1 2 3 4
M1 2 3 4 4 nmod w=100u l=10u
M2 1 2 4 4 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.ends

Va 11 0 dc 5
Vb 12 0 dc 5
Vc 13 0 dc 5
Vd 14 0 dc 0
Vdd 2 0 dc 5V
Xb 12 2 15 inverter
Xc 13 2 17 inverter
Xd 14 2 19 inverter
Xab 11 12 15 16 pass_and
Xabc 16 13 17 18 pass_and
Xabc_d 18 14 19 20 pass_or
.tran 0.1m 20m
.control
run
plot v(14)
plot V(20)
.endc
.end